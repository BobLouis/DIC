library verilog;
use verilog.vl_types.all;
entity textfixture is
end textfixture;
